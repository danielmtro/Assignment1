module game_logic_tester	(

);