module top_level(
	input 	button,
	output	led_r,
	output [6:0]  display0,
	output [6:0]  display1,
	output [6:0]  display2,
	output [6:0]  display3,
);


endmodule